`timescale 1ns / 1ps
module Pause(
	input clk, 
	output out
    );

assign out = 1'b1;

endmodule
